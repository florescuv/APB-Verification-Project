package afvip_package;

    import uvm_pkg::*;

`include "uvm_macros.svh"
`include "afvip_item.svh"
// `include "afvip_rst_item.svh"
`include "afvip_sequencer.svh"
// `include "afvip_rst_sequencer.svh"
`include "afvip_driver.svh"
// `include "afvip_rst_driver.svh"
`include "afvip_monitor.svh"
// `include "afvip_rst_monitor.svh"
// `include "afvip_passive_monitor.svh"
`include "afvip_agent.svh"
// `include "afvip_rst_agent.svh"
// `include "afvip_passive_agent_interrupt.svh"
// `include "afvip_scoreboard.svh"
// `include "afvip_environment.svh"
// `include "afvip_sequence.svh"
`include "afvip_apb_sequence_lib.svh"
// `include "afvip_rst_sequence.svh"
// `include "afvip_test.svh"
`include "afvip_coverage.svh"

    endpackage 