package afvip_tb_package;

    import uvm_pkg::*;
    `include "uvm_macros.svh"

    import afvip_package::*;
    import afvip_hw_rst_package::*;    
    import afvip_intr_package::*;
    
// `include "afvip_coverage.svh"   
`include "afvip_scoreboard.svh"
`include "afvip_environment.svh"
 
`include "afvip_virtual_sequencer.svh"

    endpackage