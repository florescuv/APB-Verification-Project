// ---------------------------------------------------------------------------------------------------------------------
// Module name: afvip_rst_interface
// HDL        : UVM
// Author     : Florescu Vlad-Andrei
// Description: It is a way to encapsulate signals into a block. All related signals are grouped together to form an interface block so that the same interface.
// Date       : 28 June, 2023
// ---------------------------------------------------------------------------------------------------------------------

interface afvip_rst_interface

(
    input clk
);

reg intf_reset;



endinterface 