package afvip_hw_rst_package;

    import uvm_pkg::*;

`include "afvip_rst_item.svh"
`include "afvip_rst_sequencer.svh"
`include "afvip_rst_driver.svh"
`include "afvip_rst_monitor.svh"
`include "afvip_rst_agent.svh"
`include "afvip_rst_sequence.svh"


endpackage 