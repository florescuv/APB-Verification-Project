package afvip_intr_package;

    import uvm_pkg::*;

`include "uvm_macros.svh"

`include "afvip_inter_item.svh"
`include "afvip_passive_monitor.svh"
`include "afvip_passive_agent_interrupt.svh"
`include "afvip_inter_coverage.svh"



    endpackage 