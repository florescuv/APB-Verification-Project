package afvip_test_package;

`include "uvm_macros.svh"
    import uvm_pkg::*;
    import afvip_package::*;
    import afvip_hw_rst_package::*;    
    import afvip_intr_package::*;
    import afvip_tb_package::*;
    
 //   `include "afvip_test.svh"
     `include "afvip_virtual_sequence.svh"
     `include "afvip_test_lib.svh"

    
endpackage 